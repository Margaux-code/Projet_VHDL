compteur_inst : compteur PORT MAP (
		clock	 => clock_sig,
		q	 => q_sig
	);
